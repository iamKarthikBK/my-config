package TB;
    module mkTb(Empty);
        Ifc_mme#(2048,128) rsa_mod <-mkMME;
        Reg#(Bool) rdy <- mkReg(False);
        rule rl_start(!rdy);
        //rsa_mod.mmeExp(1024'd211023, 1024'd101232, 1024'd410431, 1024'd25);
        let a = 2048'h3EF8F0B6A84A7C9F60C53609493A6E5D97550553669A8FF328051AD8918A29A7C714E0F32DDC5C12097C53F50EAE335EEF73081E66D54AC2334C278E016417DD9E562BFA43B11E3913B923D6162F0D9D0779D53EE54C2CC7F7A57982DE24755209FCF142CC0062DC51F0567FDD21312CCEE613EFF40597E20980E8E2E7972067D771ED20A7DFCA15727B777A243E19335404A6DBB0FBAC64D73AC9F1436E40BED14745E6DFC26C8BB7813901CB1D9FF2FFE49D72C542E7DB928DF7E46F7CBB54C60862B1FFDEA43767956F1C8F46F0952E5BAA83FCA5ADB92C9C555E1160648F97B129E1FA121B20BFAA7631E79366E8A1211364E90AA492F820D620F7ECCEB8;
        let d = 2048'h10001;
        let n = 2048'hDBC6686641E484AD414CAC014AA5735FE6BC4382438EDBDA4E0B0712E03D2E0058A64126828D0A9157B761B563469BA4388B06D4D3EF129DF72F98806C141E049D8A7AED75063BF585F6F26F04E2A6060C41FC3336FC0D6C316DBEF1DE4E16AE095F470404A15298089BCB9EFB6F71FB903374D9B2C1849BF805780278DFC49D2C801D0BB6EEDD7B3445BDF3D6F14BE26E408DBC2B65FFA9F74882929378E7F52C1837BD35AF9EF346CFB93E4ADBE96245BEBBF260416C82B2E6EC5073294D64DFAAF29084EDDCADE68BE1BBE4387F4EE0D1297B44F553EB03EBFA2589592F74ADCD29BB961AE1A32BCB00F5793F132B552CDE09A829CFF240A5F85EB30B9467;
        let rr = 2048'h5F1BAFAEF256B913445FE4514483574C86782E756C82038423AB46592E99C34E85F1A4F59070588F214AED12F0A479EBDE82ACF55CA7C29D5501691DEBC736A4E57A88B2BC6463F151C7F6F9355862AB56E258B3B161DBB6663568B19D8C70B1D2CD9AE9ADA2F0907E8C01D3C388CC73A96E0DFFB75A1F0E168D932794D27811F6B59A7531C3BAF8D68C5CA763407C3602E466BD2155BF5D77CD0360F2BDBE60949B72DF09B72AEDE8CB9F1D0FAF40929831A8E9C292E69D06576E9751EF3C228DD3C6F1BE06E716BC6E86AC483DBB8D3DA82855E8FB45653A3B8296E414F141F1C7774E2E38C1D36154A21083D99F28E0A7823CFD10F86398D35C6C55627C06;

        //let a = 128'h3EF8F0B6A84A7C9F60C53609493A6E5D;
        //let d = 128'h10001;
        //let n = 128'h4EF8F0B6A84A7C9F60C53609493A6E5D;
        //let rr = 128'd84342486036352056769109228323799158176;
        rsa_mod.mmeExp(a,d,n,rr);
        //3ef8f0b6a84a7c9f60c53609493a6e5d
        //211310595204847329841774944651329564253

        //rsa_mod.mmeExp(2048'd211023, 2048'd101232, 2048'd410431, 2048'd269910);
        //rsa_mod.mmeExp(2048'd23, 2048'd10, 2048'd101, 2048'd19);
        $display("a: %h", a);
        $display("d: %h", d);
        $display("n: %h", n);
        $display("r: %h", rr);
        rdy <= True;
        endrule

        rule rl_get_result (rdy);
        if(rsa_mod.isReady) begin
            $display($time, "Result:  %h", rsa_mod.getResult);
            $finish(0);
        end
        endrule
    endmodule
endpackage: TB