package RegArray;

    

endpackage: RegArray