package TB;

    import ModExpt :: * ;

    module mk_TB(Empty);

    endmodule: mk_TB

endpackage: TB