package junk;

import Gearbox :: *;



endpackage: junk