package tb;
endpackage: tb