package TB;

    import ModExpt :: * ;

    module mk_TB(Empty);
        ModExpt modexpt <- mkModExpt();
    endmodule: mk_TB

endpackage: TB