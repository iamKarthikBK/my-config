package ECC_template_32;
    import axi4 :: * ;
    import axi4l :: * ;
    import apb :: * ;
    import ECC :: * ;

    `define aw 32
    `define dw 32
    `define uw 0
    `define in_depth 4
    `define out_depth 5
    `define base 'h12300
endpackage: ECC_template_32