package field_ops;

    `include "acce;.defines"
    import primitives :: * ;

endpackage: field_ops