package RegV;

    import Vector :: * ;

    interface RegV;
    endinterface: RegV

endpackage: RegV