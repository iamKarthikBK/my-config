package ECC_template_32;
    import axi4 :: * ;
endpackage: ECC_template_32