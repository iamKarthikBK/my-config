package adder;

endpackage: adder