package RegArray;

    import Vector :: * ;

endpackage: RegArray